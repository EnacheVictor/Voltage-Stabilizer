** Profile: "SCHEMATIC1-sim- Vout"  [ C:\Users\Enach\Desktop\P1_2024_434D_Enache_Victor_SERS_N10_Orcad\Schematics\Proiect\proiect1_enachevictor-pspicefiles\schematic1\sim- vout.sim ] 

** Creating circuit file "sim- Vout.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../biblioteci spice/bc846b.lib" 
.LIB "../../../biblioteci spice/bc856b.lib" 
.LIB "../../../biblioteci spice/opto.lib" 
.LIB "../../../biblioteci spice/bzx84c2v7.lib" 
.LIB "../../../biblioteci spice/mjd31cg.lib" 
* From [PSPICE NETLIST] section of C:\Users\Enach\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM SET 0 1 0.01 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
